** sch_path: /home/raditya/Silicons/Projects/simple_inverter.sch
**.subckt simple_inverter
V1 VDD GND 16
V2 input GND 0
XM2 output input VDD VDD sky130_fd_pr__pfet_20v0 L=0.5 W=60 m=1
XM3 output input GND GND sky130_fd_pr__nfet_20v0_nvt W=40 L=0.5 m=1
**** begin user architecture code
 .lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt
.param mc_mmm_cwitch=0
.param mc_pr_switch=1



.option wnflag=0
.option savecurrents
.control
save all
dc v2 0 20 0.05
plot input output
op
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
