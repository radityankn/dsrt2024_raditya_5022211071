magic
tech sky130A
timestamp 1714402843
<< nwell >>
rect -95 20 60 110
rect 195 20 350 110
rect 485 20 640 110
rect 775 20 930 110
rect 1065 20 1220 110
rect -95 -195 60 -110
rect 195 -195 350 -110
rect 485 -195 640 -110
rect 775 -195 930 -110
rect 1065 -195 1220 -110
<< nmos >>
rect -20 -60 -5 -15
rect 270 -60 285 -15
rect 560 -60 575 -15
rect 850 -60 865 -15
rect 1140 -60 1155 -15
<< pmos >>
rect -20 40 -5 90
rect 270 40 285 90
rect 560 40 575 90
rect 850 40 865 90
rect 1140 40 1155 90
<< ndiff >>
rect -60 185 45 195
rect -60 155 -50 185
rect 35 155 45 185
rect -60 145 45 155
rect 230 185 335 195
rect 230 155 240 185
rect 325 155 335 185
rect 230 145 335 155
rect 520 185 625 195
rect 520 155 530 185
rect 615 155 625 185
rect 520 145 625 155
rect 810 185 915 195
rect 810 155 820 185
rect 905 155 915 185
rect 810 145 915 155
rect 1100 185 1205 195
rect 1100 155 1110 185
rect 1195 155 1205 185
rect 1100 145 1205 155
rect -65 -25 -20 -15
rect -65 -50 -55 -25
rect -35 -50 -20 -25
rect -65 -60 -20 -50
rect -5 -25 40 -15
rect -5 -50 10 -25
rect 30 -50 40 -25
rect -5 -60 40 -50
rect 225 -25 270 -15
rect 225 -50 235 -25
rect 255 -50 270 -25
rect 225 -60 270 -50
rect 285 -25 330 -15
rect 285 -50 300 -25
rect 320 -50 330 -25
rect 285 -60 330 -50
rect 515 -25 560 -15
rect 515 -50 525 -25
rect 545 -50 560 -25
rect 515 -60 560 -50
rect 575 -25 620 -15
rect 575 -50 590 -25
rect 610 -50 620 -25
rect 575 -60 620 -50
rect 805 -25 850 -15
rect 805 -50 815 -25
rect 835 -50 850 -25
rect 805 -60 850 -50
rect 865 -25 910 -15
rect 865 -50 880 -25
rect 900 -50 910 -25
rect 865 -60 910 -50
rect 1095 -25 1140 -15
rect 1095 -50 1105 -25
rect 1125 -50 1140 -25
rect 1095 -60 1140 -50
rect 1155 -25 1200 -15
rect 1155 -50 1170 -25
rect 1190 -50 1200 -25
rect 1155 -60 1200 -50
<< pdiff >>
rect -60 80 -20 90
rect -60 50 -50 80
rect -30 50 -20 80
rect -60 40 -20 50
rect -5 80 40 90
rect -5 50 10 80
rect 30 50 40 80
rect -5 40 40 50
rect 230 80 270 90
rect 230 50 240 80
rect 260 50 270 80
rect 230 40 270 50
rect 285 80 330 90
rect 285 50 300 80
rect 320 50 330 80
rect 285 40 330 50
rect 520 80 560 90
rect 520 50 530 80
rect 550 50 560 80
rect 520 40 560 50
rect 575 80 620 90
rect 575 50 590 80
rect 610 50 620 80
rect 575 40 620 50
rect 810 80 850 90
rect 810 50 820 80
rect 840 50 850 80
rect 810 40 850 50
rect 865 80 910 90
rect 865 50 880 80
rect 900 50 910 80
rect 865 40 910 50
rect 1100 80 1140 90
rect 1100 50 1110 80
rect 1130 50 1140 80
rect 1100 40 1140 50
rect 1155 80 1200 90
rect 1155 50 1170 80
rect 1190 50 1200 80
rect 1155 40 1200 50
rect -65 -135 40 -130
rect -65 -170 -55 -135
rect 30 -170 40 -135
rect -65 -175 40 -170
rect 225 -135 330 -130
rect 225 -170 235 -135
rect 320 -170 330 -135
rect 225 -175 330 -170
rect 515 -135 620 -130
rect 515 -170 525 -135
rect 610 -170 620 -135
rect 515 -175 620 -170
rect 805 -135 910 -130
rect 805 -170 815 -135
rect 900 -170 910 -135
rect 805 -175 910 -170
rect 1095 -135 1200 -130
rect 1095 -170 1105 -135
rect 1190 -170 1200 -135
rect 1095 -175 1200 -170
<< ndiffc >>
rect -50 155 35 185
rect 240 155 325 185
rect 530 155 615 185
rect 820 155 905 185
rect 1110 155 1195 185
rect -55 -50 -35 -25
rect 10 -50 30 -25
rect 235 -50 255 -25
rect 300 -50 320 -25
rect 525 -50 545 -25
rect 590 -50 610 -25
rect 815 -50 835 -25
rect 880 -50 900 -25
rect 1105 -50 1125 -25
rect 1170 -50 1190 -25
<< pdiffc >>
rect -50 50 -30 80
rect 10 50 30 80
rect 240 50 260 80
rect 300 50 320 80
rect 530 50 550 80
rect 590 50 610 80
rect 820 50 840 80
rect 880 50 900 80
rect 1110 50 1130 80
rect 1170 50 1190 80
rect -55 -170 30 -135
rect 235 -170 320 -135
rect 525 -170 610 -135
rect 815 -170 900 -135
rect 1105 -170 1190 -135
<< poly >>
rect -20 90 -5 105
rect 270 90 285 105
rect 560 90 575 105
rect 850 90 865 105
rect 1140 90 1155 105
rect -120 30 -85 35
rect -20 30 -5 40
rect 170 30 205 35
rect 270 30 285 40
rect 460 30 495 35
rect 560 30 575 40
rect 750 30 785 35
rect 850 30 865 40
rect 1040 30 1075 35
rect 1140 30 1155 40
rect -120 25 5 30
rect -120 0 -110 25
rect -90 0 5 25
rect -120 -5 5 0
rect 170 25 295 30
rect 170 0 180 25
rect 200 0 295 25
rect 170 -5 295 0
rect 460 25 585 30
rect 460 0 470 25
rect 490 0 585 25
rect 460 -5 585 0
rect 750 25 875 30
rect 750 0 760 25
rect 780 0 875 25
rect 750 -5 875 0
rect 1040 25 1165 30
rect 1040 0 1050 25
rect 1070 0 1165 25
rect 1040 -5 1165 0
rect -120 -10 -85 -5
rect -20 -15 -5 -5
rect 170 -10 205 -5
rect 270 -15 285 -5
rect 460 -10 495 -5
rect 560 -15 575 -5
rect 750 -10 785 -5
rect 850 -15 865 -5
rect 1040 -10 1075 -5
rect 1140 -15 1155 -5
rect -20 -75 -5 -60
rect 270 -75 285 -60
rect 560 -75 575 -60
rect 850 -75 865 -60
rect 1140 -75 1155 -60
<< polycont >>
rect -110 0 -90 25
rect 180 0 200 25
rect 470 0 490 25
rect 760 0 780 25
rect 1050 0 1070 25
<< locali >>
rect -60 190 45 195
rect -60 155 -50 190
rect 35 155 45 190
rect -60 145 45 155
rect 230 190 335 195
rect 230 155 240 190
rect 325 155 335 190
rect 230 145 335 155
rect 520 190 625 195
rect 520 155 530 190
rect 615 155 625 190
rect 520 145 625 155
rect 810 190 915 195
rect 810 155 820 190
rect 905 155 915 190
rect 810 145 915 155
rect 1100 190 1205 195
rect 1100 155 1110 190
rect 1195 155 1205 190
rect 1100 145 1205 155
rect -60 80 -20 145
rect -60 50 -50 80
rect -30 50 -20 80
rect -60 40 -20 50
rect 0 80 50 90
rect 0 50 10 80
rect 30 50 50 80
rect 0 40 50 50
rect 230 80 270 145
rect 230 50 240 80
rect 260 50 270 80
rect 230 40 270 50
rect 290 80 340 90
rect 290 50 300 80
rect 320 50 340 80
rect 290 40 340 50
rect 520 80 560 145
rect 520 50 530 80
rect 550 50 560 80
rect 520 40 560 50
rect 580 80 630 90
rect 580 50 590 80
rect 610 50 630 80
rect 580 40 630 50
rect 810 80 850 145
rect 810 50 820 80
rect 840 50 850 80
rect 810 40 850 50
rect 870 80 920 90
rect 870 50 880 80
rect 900 50 920 80
rect 870 40 920 50
rect 1100 80 1140 145
rect 1100 50 1110 80
rect 1130 50 1140 80
rect 1100 40 1140 50
rect 1160 80 1210 90
rect 1160 50 1170 80
rect 1190 50 1210 80
rect 1160 40 1210 50
rect 15 35 50 40
rect 305 35 340 40
rect 595 35 630 40
rect 885 35 920 40
rect 1175 35 1210 40
rect -120 30 -85 35
rect -120 -5 -115 30
rect -90 -5 -85 30
rect -120 -10 -85 -5
rect 15 -10 20 35
rect 45 -10 50 35
rect 170 30 205 35
rect 170 -5 175 30
rect 200 -5 205 30
rect 170 -10 205 -5
rect 305 -10 310 35
rect 335 -10 340 35
rect 460 30 495 35
rect 460 -5 465 30
rect 490 -5 495 30
rect 460 -10 495 -5
rect 595 -10 600 35
rect 625 -10 630 35
rect 750 30 785 35
rect 750 -5 755 30
rect 780 -5 785 30
rect 750 -10 785 -5
rect 885 -10 890 35
rect 915 -10 920 35
rect 1040 30 1075 35
rect 1040 -5 1045 30
rect 1070 -5 1075 30
rect 1040 -10 1075 -5
rect 1175 -10 1180 35
rect 1205 -10 1210 35
rect 15 -15 50 -10
rect 305 -15 340 -10
rect 595 -15 630 -10
rect 885 -15 920 -10
rect 1175 -15 1210 -10
rect -65 -25 -25 -15
rect -65 -50 -55 -25
rect -35 -50 -25 -25
rect -65 -130 -25 -50
rect 0 -25 50 -15
rect 0 -50 10 -25
rect 30 -50 50 -25
rect 0 -60 50 -50
rect 225 -25 265 -15
rect 225 -50 235 -25
rect 255 -50 265 -25
rect 225 -130 265 -50
rect 290 -25 340 -15
rect 290 -50 300 -25
rect 320 -50 340 -25
rect 290 -60 340 -50
rect 515 -25 555 -15
rect 515 -50 525 -25
rect 545 -50 555 -25
rect 515 -130 555 -50
rect 580 -25 630 -15
rect 580 -50 590 -25
rect 610 -50 630 -25
rect 580 -60 630 -50
rect 805 -25 845 -15
rect 805 -50 815 -25
rect 835 -50 845 -25
rect 805 -130 845 -50
rect 870 -25 920 -15
rect 870 -50 880 -25
rect 900 -50 920 -25
rect 870 -60 920 -50
rect 1095 -25 1135 -15
rect 1095 -50 1105 -25
rect 1125 -50 1135 -25
rect 1095 -130 1135 -50
rect 1160 -25 1210 -15
rect 1160 -50 1170 -25
rect 1190 -50 1210 -25
rect 1160 -60 1210 -50
rect -65 -135 40 -130
rect -65 -170 -55 -135
rect 30 -170 40 -135
rect -65 -175 40 -170
rect 225 -135 330 -130
rect 225 -170 235 -135
rect 320 -170 330 -135
rect 225 -175 330 -170
rect 515 -135 620 -130
rect 515 -170 525 -135
rect 610 -170 620 -135
rect 515 -175 620 -170
rect 805 -135 910 -130
rect 805 -170 815 -135
rect 900 -170 910 -135
rect 805 -175 910 -170
rect 1095 -135 1200 -130
rect 1095 -170 1105 -135
rect 1190 -170 1200 -135
rect 1095 -175 1200 -170
<< viali >>
rect -50 185 35 190
rect -50 155 35 185
rect 240 185 325 190
rect 240 155 325 185
rect 530 185 615 190
rect 530 155 615 185
rect 820 185 905 190
rect 820 155 905 185
rect 1110 185 1195 190
rect 1110 155 1195 185
rect -115 25 -90 30
rect -115 0 -110 25
rect -110 0 -90 25
rect -115 -5 -90 0
rect 20 -10 45 35
rect 175 25 200 30
rect 175 0 180 25
rect 180 0 200 25
rect 175 -5 200 0
rect 310 -10 335 35
rect 465 25 490 30
rect 465 0 470 25
rect 470 0 490 25
rect 465 -5 490 0
rect 600 -10 625 35
rect 755 25 780 30
rect 755 0 760 25
rect 760 0 780 25
rect 755 -5 780 0
rect 890 -10 915 35
rect 1045 25 1070 30
rect 1045 0 1050 25
rect 1050 0 1070 25
rect 1045 -5 1070 0
rect 1180 -10 1205 35
rect -55 -170 30 -135
rect 235 -170 320 -135
rect 525 -170 610 -135
rect 815 -170 900 -135
rect 1105 -170 1190 -135
<< metal1 >>
rect -170 190 1280 195
rect -170 155 -50 190
rect 35 155 240 190
rect 325 155 530 190
rect 615 155 820 190
rect 905 155 1110 190
rect 1195 155 1280 190
rect -170 145 1280 155
rect -170 35 -85 45
rect -170 -10 -160 35
rect -120 30 -85 35
rect -120 -5 -115 30
rect -90 -5 -85 30
rect -120 -10 -85 -5
rect -170 -20 -85 -10
rect 15 35 205 45
rect 15 -10 20 35
rect 45 30 205 35
rect 45 -5 175 30
rect 200 -5 205 30
rect 45 -10 205 -5
rect 15 -20 205 -10
rect 305 35 495 45
rect 305 -10 310 35
rect 335 30 495 35
rect 335 -5 465 30
rect 490 -5 495 30
rect 335 -10 495 -5
rect 305 -20 495 -10
rect 595 35 785 45
rect 595 -10 600 35
rect 625 30 785 35
rect 625 -5 755 30
rect 780 -5 785 30
rect 625 -10 785 -5
rect 595 -20 785 -10
rect 885 35 1075 45
rect 885 -10 890 35
rect 915 30 1075 35
rect 915 -5 1045 30
rect 1070 -5 1075 30
rect 915 -10 1075 -5
rect 885 -20 1075 -10
rect 1175 35 1345 45
rect 1175 -10 1180 35
rect 1205 -10 1230 35
rect 1270 -10 1345 35
rect 1175 -20 1345 -10
rect -170 -135 1280 -130
rect -170 -170 -55 -135
rect 30 -170 235 -135
rect 320 -170 525 -135
rect 610 -170 815 -135
rect 900 -170 1105 -135
rect 1190 -170 1280 -135
rect -170 -175 1280 -170
<< via1 >>
rect -160 -10 -120 35
rect 1230 -10 1270 35
<< metal2 >>
rect -170 35 1280 45
rect -170 -10 -160 35
rect -120 -10 1230 35
rect 1270 -10 1280 35
rect -170 -20 1280 -10
<< labels >>
rlabel metal1 80 -170 90 -160 1 vss
rlabel via1 -155 0 -145 10 1 in1
rlabel metal1 60 150 115 175 1 vdd
rlabel metal1 370 -170 380 -160 1 vss
rlabel metal1 370 5 380 15 1 out1
rlabel metal1 350 150 405 175 1 vdd
rlabel metal1 660 -170 670 -160 1 vss
rlabel metal1 660 5 670 15 1 out1
rlabel metal1 640 150 695 175 1 vdd
rlabel metal1 950 -170 960 -160 1 vss
rlabel metal1 950 5 960 15 1 out1
rlabel metal1 930 150 985 175 1 vdd
rlabel metal1 1240 -170 1250 -160 1 vss
rlabel metal1 1220 150 1275 175 1 vdd
rlabel metal1 950 5 960 15 1 out4
rlabel metal1 660 5 670 15 1 out3
rlabel metal1 370 5 380 15 1 out2
rlabel metal1 80 5 90 15 1 out1
rlabel via1 -155 0 -145 10 1 input
rlabel metal1 1325 -5 1335 5 1 output
<< end >>
