magic
tech sky130A
timestamp 1714383862
<< nwell >>
rect -85 -230 95 -145
<< nmos >>
rect -10 -110 30 -65
<< ndiff >>
rect -65 -75 -10 -65
rect -65 -95 -50 -75
rect -25 -95 -10 -75
rect -65 -110 -10 -95
rect 30 -75 80 -65
rect 30 -95 45 -75
rect 65 -95 80 -75
rect 30 -110 80 -95
<< pdiff >>
rect -65 -170 75 -165
rect -65 -190 -55 -170
rect 65 -190 75 -170
rect -65 -195 75 -190
<< ndiffc >>
rect -50 -95 -25 -75
rect 45 -95 65 -75
<< pdiffc >>
rect -55 -190 65 -170
<< poly >>
rect -10 -25 30 -20
rect -10 -45 0 -25
rect 20 -45 30 -25
rect -10 -65 30 -45
rect -10 -125 30 -110
<< polycont >>
rect 0 -45 20 -25
<< locali >>
rect -10 -25 30 -20
rect -10 -45 0 -25
rect 25 -45 30 -25
rect -10 -50 30 -45
rect -60 -75 -15 -70
rect 35 -75 75 -70
rect -60 -165 -15 -105
rect -65 -170 75 -165
rect -65 -190 -55 -170
rect 65 -190 75 -170
rect -65 -195 75 -190
<< viali >>
rect 0 -45 20 -25
rect 20 -45 25 -25
rect -60 -95 -50 -75
rect -50 -95 -25 -75
rect -25 -95 -15 -75
rect -60 -105 -15 -95
rect 35 -95 45 -75
rect 45 -95 65 -75
rect 65 -95 75 -75
rect 35 -105 75 -95
<< metal1 >>
rect -10 -25 160 -20
rect -10 -45 0 -25
rect 25 -45 160 -25
rect -10 -50 160 -45
rect -65 -75 -10 -65
rect -65 -105 -60 -75
rect -15 -105 -10 -75
rect -65 -300 -10 -105
rect 30 -75 80 -65
rect 30 -105 35 -75
rect 75 -105 80 -75
rect 30 -300 80 -105
rect 110 -300 160 -50
<< labels >>
rlabel metal1 -50 -265 -50 -265 1 gnd
rlabel metal1 45 -275 45 -275 1 vcc
rlabel metal1 140 -195 140 -195 1 in
<< end >>
